library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sid_coeffs is
  port (
    clka   : in  std_logic;
    clkb   : in  std_logic;
    addra  : in  unsigned(11 downto 0);
    addrb  : in  unsigned(11 downto 0);
    dia    : in  unsigned(7 downto 0) := (others => '0');
    dib    : in  unsigned(7 downto 0) := (others => '0');
    douta  : out unsigned(7 downto 0) := (others => 'Z');
    doutb  : out unsigned(7 downto 0) := (others => '0');
    wea    : in  std_logic;
    web    : in  std_logic;
    ena    : in  std_logic;
    enb    : in  std_logic
    -- rsta   : in  std_logic;
    -- rstb   : in  std_logic;
    -- regcea : in  std_logic;
    -- regceb : in  std_logic
    );
end entity;

architecture beh of sid_coeffs is

  type mtype is array(natural range 0 to 4095) of unsigned(7 downto 0);

  constant coef_init : mtype := (
    x"1E", x"00", x"23", x"00", x"29", x"00", x"2F", x"00", x"35", x"00", x"3B", x"00", x"41", x"00", x"46", x"00", 
    x"4C", x"00", x"52", x"00", x"58", x"00", x"5E", x"00", x"64", x"00", x"6A", x"00", x"6F", x"00", x"75", x"00", 
    x"7B", x"00", x"81", x"00", x"87", x"00", x"8D", x"00", x"92", x"00", x"98", x"00", x"9E", x"00", x"A4", x"00", 
    x"AA", x"00", x"B0", x"00", x"B6", x"00", x"BB", x"00", x"C1", x"00", x"C7", x"00", x"CD", x"00", x"D3", x"00", 
    x"D9", x"00", x"DE", x"00", x"E4", x"00", x"EA", x"00", x"F0", x"00", x"F6", x"00", x"FC", x"00", x"02", x"01", 
    x"07", x"01", x"0D", x"01", x"13", x"01", x"19", x"01", x"1F", x"01", x"25", x"01", x"2A", x"01", x"30", x"01", 
    x"36", x"01", x"3C", x"01", x"42", x"01", x"48", x"01", x"4E", x"01", x"53", x"01", x"59", x"01", x"5F", x"01", 
    x"65", x"01", x"6B", x"01", x"71", x"01", x"77", x"01", x"7C", x"01", x"82", x"01", x"88", x"01", x"8E", x"01", 
    x"94", x"01", x"9A", x"01", x"9F", x"01", x"A5", x"01", x"AB", x"01", x"B1", x"01", x"B7", x"01", x"BD", x"01", 
    x"C3", x"01", x"C8", x"01", x"CE", x"01", x"D4", x"01", x"DA", x"01", x"E0", x"01", x"E6", x"01", x"EB", x"01", 
    x"F1", x"01", x"F7", x"01", x"FD", x"01", x"03", x"02", x"09", x"02", x"0F", x"02", x"14", x"02", x"1A", x"02", 
    x"20", x"02", x"26", x"02", x"2C", x"02", x"32", x"02", x"37", x"02", x"3D", x"02", x"43", x"02", x"49", x"02", 
    x"4F", x"02", x"55", x"02", x"5B", x"02", x"60", x"02", x"66", x"02", x"6C", x"02", x"72", x"02", x"78", x"02", 
    x"7E", x"02", x"83", x"02", x"89", x"02", x"8F", x"02", x"95", x"02", x"9B", x"02", x"A1", x"02", x"A7", x"02", 
    x"AC", x"02", x"B2", x"02", x"B8", x"02", x"BE", x"02", x"C4", x"02", x"CA", x"02", x"D0", x"02", x"D5", x"02", 
    x"DB", x"02", x"E1", x"02", x"E7", x"02", x"ED", x"02", x"F3", x"02", x"F8", x"02", x"FE", x"02", x"04", x"03", 
    x"0A", x"03", x"10", x"03", x"16", x"03", x"1C", x"03", x"21", x"03", x"27", x"03", x"2D", x"03", x"33", x"03", 
    x"39", x"03", x"3F", x"03", x"44", x"03", x"4A", x"03", x"50", x"03", x"56", x"03", x"5C", x"03", x"62", x"03", 
    x"68", x"03", x"6D", x"03", x"73", x"03", x"79", x"03", x"7F", x"03", x"85", x"03", x"8B", x"03", x"90", x"03", 
    x"96", x"03", x"9C", x"03", x"A2", x"03", x"A8", x"03", x"AE", x"03", x"B4", x"03", x"B9", x"03", x"BF", x"03", 
    x"C5", x"03", x"CB", x"03", x"D1", x"03", x"D7", x"03", x"DD", x"03", x"E2", x"03", x"E8", x"03", x"EE", x"03", 
    x"F4", x"03", x"FA", x"03", x"00", x"04", x"05", x"04", x"0B", x"04", x"11", x"04", x"17", x"04", x"1D", x"04", 
    x"23", x"04", x"29", x"04", x"2E", x"04", x"34", x"04", x"3A", x"04", x"40", x"04", x"46", x"04", x"4C", x"04", 
    x"51", x"04", x"57", x"04", x"5D", x"04", x"63", x"04", x"69", x"04", x"6F", x"04", x"75", x"04", x"7A", x"04", 
    x"80", x"04", x"86", x"04", x"8C", x"04", x"92", x"04", x"98", x"04", x"9D", x"04", x"A3", x"04", x"A9", x"04", 
    x"AF", x"04", x"B5", x"04", x"BB", x"04", x"C1", x"04", x"C6", x"04", x"CC", x"04", x"D2", x"04", x"D8", x"04", 
    x"DE", x"04", x"E4", x"04", x"E9", x"04", x"EF", x"04", x"F5", x"04", x"FB", x"04", x"01", x"05", x"07", x"05", 
    x"0D", x"05", x"12", x"05", x"18", x"05", x"1E", x"05", x"24", x"05", x"2A", x"05", x"30", x"05", x"36", x"05", 
    x"3B", x"05", x"41", x"05", x"47", x"05", x"4D", x"05", x"53", x"05", x"59", x"05", x"5E", x"05", x"64", x"05", 
    x"6A", x"05", x"70", x"05", x"76", x"05", x"7C", x"05", x"82", x"05", x"87", x"05", x"8D", x"05", x"93", x"05", 
    x"99", x"05", x"9F", x"05", x"A5", x"05", x"AA", x"05", x"B0", x"05", x"B6", x"05", x"BC", x"05", x"C2", x"05", 
    x"C8", x"05", x"CE", x"05", x"D3", x"05", x"D9", x"05", x"DF", x"05", x"E5", x"05", x"EB", x"05", x"F1", x"05", 
    x"F6", x"05", x"FC", x"05", x"02", x"06", x"08", x"06", x"0E", x"06", x"14", x"06", x"1A", x"06", x"1F", x"06", 
    x"25", x"06", x"2B", x"06", x"31", x"06", x"37", x"06", x"3D", x"06", x"42", x"06", x"48", x"06", x"4E", x"06", 
    x"54", x"06", x"5A", x"06", x"60", x"06", x"66", x"06", x"6B", x"06", x"71", x"06", x"77", x"06", x"7D", x"06", 
    x"83", x"06", x"89", x"06", x"8F", x"06", x"94", x"06", x"9A", x"06", x"A0", x"06", x"A6", x"06", x"AC", x"06", 
    x"B2", x"06", x"B7", x"06", x"BD", x"06", x"C3", x"06", x"C9", x"06", x"CF", x"06", x"D5", x"06", x"DB", x"06", 
    x"E0", x"06", x"E6", x"06", x"EC", x"06", x"F2", x"06", x"F8", x"06", x"FE", x"06", x"03", x"07", x"09", x"07", 
    x"0F", x"07", x"15", x"07", x"1B", x"07", x"21", x"07", x"27", x"07", x"2C", x"07", x"32", x"07", x"38", x"07", 
    x"3E", x"07", x"44", x"07", x"4A", x"07", x"4F", x"07", x"55", x"07", x"5B", x"07", x"61", x"07", x"67", x"07", 
    x"6D", x"07", x"73", x"07", x"78", x"07", x"7E", x"07", x"84", x"07", x"8A", x"07", x"90", x"07", x"96", x"07", 
    x"9C", x"07", x"A1", x"07", x"A7", x"07", x"AD", x"07", x"B3", x"07", x"B9", x"07", x"BF", x"07", x"C4", x"07", 
    x"CA", x"07", x"D0", x"07", x"D6", x"07", x"DC", x"07", x"E2", x"07", x"E8", x"07", x"ED", x"07", x"F3", x"07", 
    x"F9", x"07", x"FF", x"07", x"05", x"08", x"0B", x"08", x"10", x"08", x"16", x"08", x"1C", x"08", x"22", x"08", 
    x"28", x"08", x"2E", x"08", x"34", x"08", x"39", x"08", x"3F", x"08", x"45", x"08", x"4B", x"08", x"51", x"08", 
    x"57", x"08", x"5C", x"08", x"62", x"08", x"68", x"08", x"6E", x"08", x"74", x"08", x"7A", x"08", x"80", x"08", 
    x"85", x"08", x"8B", x"08", x"91", x"08", x"97", x"08", x"9D", x"08", x"A3", x"08", x"A8", x"08", x"AE", x"08", 
    x"B4", x"08", x"BA", x"08", x"C0", x"08", x"C6", x"08", x"CC", x"08", x"D1", x"08", x"D7", x"08", x"DD", x"08", 
    x"E3", x"08", x"E9", x"08", x"EF", x"08", x"F5", x"08", x"FA", x"08", x"00", x"09", x"06", x"09", x"0C", x"09", 
    x"12", x"09", x"18", x"09", x"1D", x"09", x"23", x"09", x"29", x"09", x"2F", x"09", x"35", x"09", x"3B", x"09", 
    x"41", x"09", x"46", x"09", x"4C", x"09", x"52", x"09", x"58", x"09", x"5E", x"09", x"64", x"09", x"69", x"09", 
    x"6F", x"09", x"75", x"09", x"7B", x"09", x"81", x"09", x"87", x"09", x"8D", x"09", x"92", x"09", x"98", x"09", 
    x"9E", x"09", x"A4", x"09", x"AA", x"09", x"B0", x"09", x"B5", x"09", x"BB", x"09", x"C1", x"09", x"C7", x"09", 
    x"CD", x"09", x"D3", x"09", x"D9", x"09", x"DE", x"09", x"E4", x"09", x"EA", x"09", x"F0", x"09", x"F6", x"09", 
    x"FC", x"09", x"02", x"0A", x"07", x"0A", x"0D", x"0A", x"13", x"0A", x"19", x"0A", x"1F", x"0A", x"25", x"0A", 
    x"2A", x"0A", x"30", x"0A", x"36", x"0A", x"3C", x"0A", x"42", x"0A", x"48", x"0A", x"4E", x"0A", x"53", x"0A", 
    x"59", x"0A", x"5F", x"0A", x"65", x"0A", x"6B", x"0A", x"71", x"0A", x"76", x"0A", x"7C", x"0A", x"82", x"0A", 
    x"88", x"0A", x"8E", x"0A", x"94", x"0A", x"9A", x"0A", x"9F", x"0A", x"A5", x"0A", x"AB", x"0A", x"B1", x"0A", 
    x"B7", x"0A", x"BD", x"0A", x"C2", x"0A", x"C8", x"0A", x"CE", x"0A", x"D4", x"0A", x"DA", x"0A", x"E0", x"0A", 
    x"E6", x"0A", x"EB", x"0A", x"F1", x"0A", x"F7", x"0A", x"FD", x"0A", x"03", x"0B", x"09", x"0B", x"0E", x"0B", 
    x"14", x"0B", x"1A", x"0B", x"20", x"0B", x"26", x"0B", x"2C", x"0B", x"32", x"0B", x"37", x"0B", x"3D", x"0B", 
    x"43", x"0B", x"49", x"0B", x"4F", x"0B", x"55", x"0B", x"5B", x"0B", x"60", x"0B", x"66", x"0B", x"6C", x"0B", 
    x"72", x"0B", x"78", x"0B", x"7E", x"0B", x"83", x"0B", x"89", x"0B", x"8F", x"0B", x"95", x"0B", x"9B", x"0B", 
    x"A1", x"0B", x"A7", x"0B", x"AC", x"0B", x"B2", x"0B", x"B8", x"0B", x"BE", x"0B", x"C4", x"0B", x"CA", x"0B", 
    x"CF", x"0B", x"D5", x"0B", x"DB", x"0B", x"E1", x"0B", x"E7", x"0B", x"ED", x"0B", x"F3", x"0B", x"F8", x"0B", 
    x"FE", x"0B", x"04", x"0C", x"0A", x"0C", x"10", x"0C", x"16", x"0C", x"1B", x"0C", x"21", x"0C", x"27", x"0C", 
    x"2D", x"0C", x"33", x"0C", x"39", x"0C", x"3F", x"0C", x"44", x"0C", x"4A", x"0C", x"50", x"0C", x"56", x"0C", 
    x"5C", x"0C", x"62", x"0C", x"67", x"0C", x"6D", x"0C", x"73", x"0C", x"79", x"0C", x"7F", x"0C", x"85", x"0C", 
    x"8B", x"0C", x"90", x"0C", x"96", x"0C", x"9C", x"0C", x"A2", x"0C", x"A8", x"0C", x"AE", x"0C", x"B4", x"0C", 
    x"B9", x"0C", x"BF", x"0C", x"C5", x"0C", x"CB", x"0C", x"D1", x"0C", x"D7", x"0C", x"DC", x"0C", x"E2", x"0C", 
    x"E8", x"0C", x"EE", x"0C", x"F4", x"0C", x"FA", x"0C", x"00", x"0D", x"05", x"0D", x"0B", x"0D", x"11", x"0D", 
    x"17", x"0D", x"1D", x"0D", x"23", x"0D", x"28", x"0D", x"2E", x"0D", x"34", x"0D", x"3A", x"0D", x"40", x"0D", 
    x"46", x"0D", x"4C", x"0D", x"51", x"0D", x"57", x"0D", x"5D", x"0D", x"63", x"0D", x"69", x"0D", x"6F", x"0D", 
    x"74", x"0D", x"7A", x"0D", x"80", x"0D", x"86", x"0D", x"8C", x"0D", x"92", x"0D", x"98", x"0D", x"9D", x"0D", 
    x"A3", x"0D", x"A9", x"0D", x"AF", x"0D", x"B5", x"0D", x"BB", x"0D", x"C1", x"0D", x"C6", x"0D", x"CC", x"0D", 
    x"D2", x"0D", x"D8", x"0D", x"DE", x"0D", x"E4", x"0D", x"E9", x"0D", x"EF", x"0D", x"F5", x"0D", x"FB", x"0D", 
    x"01", x"0E", x"07", x"0E", x"0D", x"0E", x"12", x"0E", x"18", x"0E", x"1E", x"0E", x"24", x"0E", x"2A", x"0E", 
    x"30", x"0E", x"35", x"0E", x"3B", x"0E", x"41", x"0E", x"47", x"0E", x"4D", x"0E", x"53", x"0E", x"59", x"0E", 
    x"5E", x"0E", x"64", x"0E", x"6A", x"0E", x"70", x"0E", x"76", x"0E", x"7C", x"0E", x"81", x"0E", x"87", x"0E", 
    x"8D", x"0E", x"93", x"0E", x"99", x"0E", x"9F", x"0E", x"A5", x"0E", x"AA", x"0E", x"B0", x"0E", x"B6", x"0E", 
    x"BC", x"0E", x"C2", x"0E", x"C8", x"0E", x"CD", x"0E", x"D3", x"0E", x"D9", x"0E", x"DF", x"0E", x"E5", x"0E", 
    x"EB", x"0E", x"F1", x"0E", x"F6", x"0E", x"FC", x"0E", x"02", x"0F", x"08", x"0F", x"0E", x"0F", x"14", x"0F", 
    x"1A", x"0F", x"1F", x"0F", x"25", x"0F", x"2B", x"0F", x"31", x"0F", x"37", x"0F", x"3D", x"0F", x"42", x"0F", 
    x"48", x"0F", x"4E", x"0F", x"54", x"0F", x"5A", x"0F", x"60", x"0F", x"66", x"0F", x"6B", x"0F", x"71", x"0F", 
    x"77", x"0F", x"7D", x"0F", x"83", x"0F", x"89", x"0F", x"8E", x"0F", x"94", x"0F", x"9A", x"0F", x"A0", x"0F", 
    x"A6", x"0F", x"AC", x"0F", x"B2", x"0F", x"B7", x"0F", x"BD", x"0F", x"C3", x"0F", x"C9", x"0F", x"CF", x"0F", 
    x"D5", x"0F", x"DA", x"0F", x"E0", x"0F", x"E6", x"0F", x"EC", x"0F", x"F2", x"0F", x"F8", x"0F", x"FE", x"0F", 
    x"03", x"10", x"09", x"10", x"0F", x"10", x"15", x"10", x"1B", x"10", x"21", x"10", x"27", x"10", x"2C", x"10", 
    x"32", x"10", x"38", x"10", x"3E", x"10", x"44", x"10", x"4A", x"10", x"4F", x"10", x"55", x"10", x"5B", x"10", 
    x"61", x"10", x"67", x"10", x"6D", x"10", x"73", x"10", x"78", x"10", x"7E", x"10", x"84", x"10", x"8A", x"10", 
    x"90", x"10", x"96", x"10", x"9B", x"10", x"A1", x"10", x"A7", x"10", x"AD", x"10", x"B3", x"10", x"B9", x"10", 
    x"BF", x"10", x"C4", x"10", x"CA", x"10", x"D0", x"10", x"D6", x"10", x"DC", x"10", x"E2", x"10", x"E7", x"10", 
    x"ED", x"10", x"F3", x"10", x"F9", x"10", x"FF", x"10", x"05", x"11", x"0B", x"11", x"10", x"11", x"16", x"11", 
    x"1C", x"11", x"22", x"11", x"28", x"11", x"2E", x"11", x"33", x"11", x"39", x"11", x"3F", x"11", x"45", x"11", 
    x"4B", x"11", x"51", x"11", x"57", x"11", x"5C", x"11", x"62", x"11", x"68", x"11", x"6E", x"11", x"74", x"11", 
    x"7A", x"11", x"80", x"11", x"85", x"11", x"8B", x"11", x"91", x"11", x"97", x"11", x"9D", x"11", x"A3", x"11", 
    x"A8", x"11", x"AE", x"11", x"B4", x"11", x"BA", x"11", x"C0", x"11", x"C6", x"11", x"CC", x"11", x"D1", x"11", 
    x"D7", x"11", x"DD", x"11", x"E3", x"11", x"E9", x"11", x"EF", x"11", x"F4", x"11", x"FA", x"11", x"00", x"12", 
    x"06", x"12", x"0C", x"12", x"12", x"12", x"18", x"12", x"1D", x"12", x"23", x"12", x"29", x"12", x"2F", x"12", 
    x"35", x"12", x"3B", x"12", x"40", x"12", x"46", x"12", x"4C", x"12", x"52", x"12", x"58", x"12", x"5E", x"12", 
    x"64", x"12", x"69", x"12", x"6F", x"12", x"75", x"12", x"7B", x"12", x"81", x"12", x"87", x"12", x"8C", x"12", 
    x"92", x"12", x"98", x"12", x"9E", x"12", x"A4", x"12", x"AA", x"12", x"B0", x"12", x"B5", x"12", x"BB", x"12", 
    x"C1", x"12", x"C7", x"12", x"CD", x"12", x"D3", x"12", x"D9", x"12", x"DE", x"12", x"E4", x"12", x"EA", x"12", 
    x"F0", x"12", x"F6", x"12", x"FC", x"12", x"01", x"13", x"07", x"13", x"0D", x"13", x"13", x"13", x"19", x"13", 
    x"1F", x"13", x"25", x"13", x"2A", x"13", x"30", x"13", x"36", x"13", x"3C", x"13", x"42", x"13", x"48", x"13", 
    x"4D", x"13", x"53", x"13", x"59", x"13", x"5F", x"13", x"65", x"13", x"6B", x"13", x"71", x"13", x"76", x"13", 
    x"7C", x"13", x"82", x"13", x"88", x"13", x"8E", x"13", x"94", x"13", x"99", x"13", x"9F", x"13", x"A5", x"13", 
    x"AB", x"13", x"B1", x"13", x"B7", x"13", x"BD", x"13", x"C2", x"13", x"C8", x"13", x"CE", x"13", x"D4", x"13", 
    x"DA", x"13", x"E0", x"13", x"E6", x"13", x"EB", x"13", x"F1", x"13", x"F7", x"13", x"FD", x"13", x"03", x"14", 
    x"09", x"14", x"0E", x"14", x"14", x"14", x"1A", x"14", x"20", x"14", x"26", x"14", x"2C", x"14", x"32", x"14", 
    x"37", x"14", x"3D", x"14", x"43", x"14", x"49", x"14", x"4F", x"14", x"55", x"14", x"5A", x"14", x"60", x"14", 
    x"66", x"14", x"6C", x"14", x"72", x"14", x"78", x"14", x"7E", x"14", x"83", x"14", x"89", x"14", x"8F", x"14", 
    x"95", x"14", x"9B", x"14", x"A1", x"14", x"A6", x"14", x"AC", x"14", x"B2", x"14", x"B8", x"14", x"BE", x"14", 
    x"C4", x"14", x"CA", x"14", x"CF", x"14", x"D5", x"14", x"DB", x"14", x"E1", x"14", x"E7", x"14", x"ED", x"14", 
    x"F2", x"14", x"F8", x"14", x"FE", x"14", x"04", x"15", x"0A", x"15", x"10", x"15", x"16", x"15", x"1B", x"15", 
    x"21", x"15", x"27", x"15", x"2D", x"15", x"33", x"15", x"39", x"15", x"3F", x"15", x"44", x"15", x"4A", x"15", 
    x"50", x"15", x"56", x"15", x"5C", x"15", x"62", x"15", x"67", x"15", x"6D", x"15", x"73", x"15", x"79", x"15", 
    x"7F", x"15", x"85", x"15", x"8B", x"15", x"90", x"15", x"96", x"15", x"9C", x"15", x"A2", x"15", x"A8", x"15", 
    x"AE", x"15", x"B3", x"15", x"B9", x"15", x"BF", x"15", x"C5", x"15", x"CB", x"15", x"D1", x"15", x"D7", x"15", 
    x"DC", x"15", x"E2", x"15", x"E8", x"15", x"EE", x"15", x"F4", x"15", x"FA", x"15", x"FF", x"15", x"05", x"16", 
    x"0B", x"16", x"11", x"16", x"17", x"16", x"1D", x"16", x"23", x"16", x"28", x"16", x"2E", x"16", x"34", x"16", 
    x"3A", x"16", x"40", x"16", x"46", x"16", x"4C", x"16", x"51", x"16", x"57", x"16", x"5D", x"16", x"63", x"16", 
    x"69", x"16", x"6F", x"16", x"74", x"16", x"7A", x"16", x"80", x"16", x"86", x"16", x"8C", x"16", x"92", x"16", 
    x"98", x"16", x"9D", x"16", x"A3", x"16", x"A9", x"16", x"AF", x"16", x"B5", x"16", x"BB", x"16", x"C0", x"16", 
    x"C6", x"16", x"CC", x"16", x"D2", x"16", x"D8", x"16", x"DE", x"16", x"E4", x"16", x"E9", x"16", x"EF", x"16", 
    x"F5", x"16", x"FB", x"16", x"01", x"17", x"07", x"17", x"0C", x"17", x"12", x"17", x"18", x"17", x"1E", x"17", 
    x"24", x"17", x"2A", x"17", x"30", x"17", x"35", x"17", x"3B", x"17", x"41", x"17", x"47", x"17", x"4D", x"17", 
    x"53", x"17", x"58", x"17", x"5E", x"17", x"64", x"17", x"6A", x"17", x"70", x"17", x"76", x"17", x"7C", x"17", 
    x"81", x"17", x"87", x"17", x"8D", x"17", x"93", x"17", x"99", x"17", x"9F", x"17", x"A5", x"17", x"AA", x"17", 
    x"B0", x"17", x"B6", x"17", x"BC", x"17", x"C2", x"17", x"C8", x"17", x"CD", x"17", x"D3", x"17", x"D9", x"17", 
    x"DF", x"17", x"E5", x"17", x"EB", x"17", x"F1", x"17", x"F6", x"17", x"FC", x"17", x"02", x"18", x"08", x"18", 
    x"0E", x"18", x"14", x"18", x"19", x"18", x"1F", x"18", x"25", x"18", x"2B", x"18", x"31", x"18", x"37", x"18", 
    x"3D", x"18", x"42", x"18", x"48", x"18", x"4E", x"18", x"54", x"18", x"5A", x"18", x"60", x"18", x"65", x"18", 
    x"6B", x"18", x"71", x"18", x"77", x"18", x"7D", x"18", x"83", x"18", x"89", x"18", x"8E", x"18", x"94", x"18", 
    x"9A", x"18", x"A0", x"18", x"A6", x"18", x"AC", x"18", x"B1", x"18", x"B7", x"18", x"BD", x"18", x"C3", x"18", 
    x"C9", x"18", x"CF", x"18", x"D5", x"18", x"DA", x"18", x"E0", x"18", x"E6", x"18", x"EC", x"18", x"F2", x"18", 
    x"F8", x"18", x"FE", x"18", x"03", x"19", x"09", x"19", x"0F", x"19", x"15", x"19", x"1B", x"19", x"21", x"19", 
    x"26", x"19", x"2C", x"19", x"32", x"19", x"38", x"19", x"3E", x"19", x"44", x"19", x"4A", x"19", x"4F", x"19", 
    x"55", x"19", x"5B", x"19", x"61", x"19", x"67", x"19", x"6D", x"19", x"72", x"19", x"78", x"19", x"7E", x"19", 
    x"84", x"19", x"8A", x"19", x"90", x"19", x"96", x"19", x"9B", x"19", x"A1", x"19", x"A7", x"19", x"AD", x"19", 
    x"B3", x"19", x"B9", x"19", x"BE", x"19", x"C4", x"19", x"CA", x"19", x"D0", x"19", x"D6", x"19", x"DC", x"19", 
    x"E2", x"19", x"E7", x"19", x"ED", x"19", x"F3", x"19", x"F9", x"19", x"FF", x"19", x"05", x"1A", x"0B", x"1A", 
    x"10", x"1A", x"16", x"1A", x"1C", x"1A", x"22", x"1A", x"28", x"1A", x"2E", x"1A", x"33", x"1A", x"39", x"1A", 
    x"3F", x"1A", x"45", x"1A", x"4B", x"1A", x"51", x"1A", x"57", x"1A", x"5C", x"1A", x"62", x"1A", x"68", x"1A", 
    x"6E", x"1A", x"74", x"1A", x"7A", x"1A", x"7F", x"1A", x"85", x"1A", x"8B", x"1A", x"91", x"1A", x"97", x"1A", 
    x"9D", x"1A", x"A3", x"1A", x"A8", x"1A", x"AE", x"1A", x"B4", x"1A", x"BA", x"1A", x"C0", x"1A", x"C6", x"1A", 
    x"CB", x"1A", x"D1", x"1A", x"D7", x"1A", x"DD", x"1A", x"E3", x"1A", x"E9", x"1A", x"EF", x"1A", x"F4", x"1A", 
    x"FA", x"1A", x"00", x"1B", x"06", x"1B", x"0C", x"1B", x"12", x"1B", x"17", x"1B", x"1D", x"1B", x"23", x"1B", 
    x"29", x"1B", x"2F", x"1B", x"35", x"1B", x"3B", x"1B", x"40", x"1B", x"46", x"1B", x"4C", x"1B", x"52", x"1B", 
    x"58", x"1B", x"5E", x"1B", x"64", x"1B", x"69", x"1B", x"6F", x"1B", x"75", x"1B", x"7B", x"1B", x"81", x"1B", 
    x"87", x"1B", x"8C", x"1B", x"92", x"1B", x"98", x"1B", x"9E", x"1B", x"A4", x"1B", x"AA", x"1B", x"B0", x"1B", 
    x"B5", x"1B", x"BB", x"1B", x"C1", x"1B", x"C7", x"1B", x"CD", x"1B", x"D3", x"1B", x"D8", x"1B", x"DE", x"1B", 
    x"E4", x"1B", x"EA", x"1B", x"F0", x"1B", x"F6", x"1B", x"FC", x"1B", x"01", x"1C", x"07", x"1C", x"0D", x"1C", 
    x"13", x"1C", x"19", x"1C", x"1F", x"1C", x"24", x"1C", x"2A", x"1C", x"30", x"1C", x"36", x"1C", x"3C", x"1C", 
    x"42", x"1C", x"48", x"1C", x"4D", x"1C", x"53", x"1C", x"59", x"1C", x"5F", x"1C", x"65", x"1C", x"6B", x"1C", 
    x"71", x"1C", x"76", x"1C", x"7C", x"1C", x"82", x"1C", x"88", x"1C", x"8E", x"1C", x"94", x"1C", x"99", x"1C", 
    x"9F", x"1C", x"A5", x"1C", x"AB", x"1C", x"B1", x"1C", x"B7", x"1C", x"BD", x"1C", x"C2", x"1C", x"C8", x"1C", 
    x"CE", x"1C", x"D4", x"1C", x"DA", x"1C", x"E0", x"1C", x"E5", x"1C", x"EB", x"1C", x"F1", x"1C", x"F7", x"1C", 
    x"FD", x"1C", x"03", x"1D", x"09", x"1D", x"0E", x"1D", x"14", x"1D", x"1A", x"1D", x"20", x"1D", x"26", x"1D", 
    x"2C", x"1D", x"31", x"1D", x"37", x"1D", x"3D", x"1D", x"43", x"1D", x"49", x"1D", x"4F", x"1D", x"55", x"1D", 
    x"5A", x"1D", x"60", x"1D", x"66", x"1D", x"6C", x"1D", x"72", x"1D", x"78", x"1D", x"7D", x"1D", x"83", x"1D", 
    x"89", x"1D", x"8F", x"1D", x"95", x"1D", x"9B", x"1D", x"A1", x"1D", x"A6", x"1D", x"AC", x"1D", x"B2", x"1D", 
    x"B8", x"1D", x"BE", x"1D", x"C4", x"1D", x"CA", x"1D", x"CF", x"1D", x"D5", x"1D", x"DB", x"1D", x"E1", x"1D", 
    x"E7", x"1D", x"ED", x"1D", x"F2", x"1D", x"F8", x"1D", x"FE", x"1D", x"04", x"1E", x"0A", x"1E", x"10", x"1E", 
    x"16", x"1E", x"1B", x"1E", x"21", x"1E", x"27", x"1E", x"2D", x"1E", x"33", x"1E", x"39", x"1E", x"3E", x"1E", 
    x"44", x"1E", x"4A", x"1E", x"50", x"1E", x"56", x"1E", x"5C", x"1E", x"62", x"1E", x"67", x"1E", x"6D", x"1E", 
    x"73", x"1E", x"79", x"1E", x"7F", x"1E", x"85", x"1E", x"8A", x"1E", x"90", x"1E", x"96", x"1E", x"9C", x"1E", 
    x"A2", x"1E", x"A8", x"1E", x"AE", x"1E", x"B3", x"1E", x"B9", x"1E", x"BF", x"1E", x"C5", x"1E", x"CB", x"1E", 
    x"D1", x"1E", x"D6", x"1E", x"DC", x"1E", x"E2", x"1E", x"E8", x"1E", x"EE", x"1E", x"F4", x"1E", x"FA", x"1E", 
    x"FF", x"1E", x"05", x"1F", x"0B", x"1F", x"11", x"1F", x"17", x"1F", x"1D", x"1F", x"23", x"1F", x"28", x"1F", 
    x"2E", x"1F", x"34", x"1F", x"3A", x"1F", x"40", x"1F", x"46", x"1F", x"4B", x"1F", x"51", x"1F", x"57", x"1F", 
    x"5D", x"1F", x"63", x"1F", x"69", x"1F", x"6F", x"1F", x"74", x"1F", x"7A", x"1F", x"80", x"1F", x"86", x"1F", 
    x"8C", x"1F", x"92", x"1F", x"97", x"1F", x"9D", x"1F", x"A3", x"1F", x"A9", x"1F", x"AF", x"1F", x"B5", x"1F", 
    x"BB", x"1F", x"C0", x"1F", x"C6", x"1F", x"CC", x"1F", x"D2", x"1F", x"D8", x"1F", x"DE", x"1F", x"E3", x"1F", 
    x"E9", x"1F", x"EF", x"1F", x"F5", x"1F", x"FB", x"1F", x"01", x"20", x"07", x"20", x"0C", x"20", x"12", x"20", 
    x"18", x"20", x"1E", x"20", x"24", x"20", x"2A", x"20", x"30", x"20", x"35", x"20", x"3B", x"20", x"41", x"20", 
    x"47", x"20", x"4D", x"20", x"53", x"20", x"58", x"20", x"5E", x"20", x"64", x"20", x"6A", x"20", x"70", x"20", 
    x"76", x"20", x"7C", x"20", x"81", x"20", x"87", x"20", x"8D", x"20", x"93", x"20", x"99", x"20", x"9F", x"20", 
    x"A4", x"20", x"AA", x"20", x"B0", x"20", x"B6", x"20", x"BC", x"20", x"C2", x"20", x"C8", x"20", x"CD", x"20", 
    x"D3", x"20", x"D9", x"20", x"DF", x"20", x"E5", x"20", x"EB", x"20", x"F0", x"20", x"F6", x"20", x"FC", x"20", 
    x"02", x"21", x"08", x"21", x"0E", x"21", x"14", x"21", x"19", x"21", x"1F", x"21", x"25", x"21", x"2B", x"21", 
    x"31", x"21", x"37", x"21", x"3C", x"21", x"42", x"21", x"48", x"21", x"4E", x"21", x"54", x"21", x"5A", x"21", 
    x"60", x"21", x"65", x"21", x"6B", x"21", x"71", x"21", x"77", x"21", x"7D", x"21", x"83", x"21", x"89", x"21", 
    x"8E", x"21", x"94", x"21", x"9A", x"21", x"A0", x"21", x"A6", x"21", x"AC", x"21", x"B1", x"21", x"B7", x"21", 
    x"BD", x"21", x"C3", x"21", x"C9", x"21", x"CF", x"21", x"D5", x"21", x"DA", x"21", x"E0", x"21", x"E6", x"21", 
    x"EC", x"21", x"F2", x"21", x"F8", x"21", x"FD", x"21", x"03", x"22", x"09", x"22", x"0F", x"22", x"15", x"22", 
    x"1B", x"22", x"21", x"22", x"26", x"22", x"2C", x"22", x"32", x"22", x"38", x"22", x"3E", x"22", x"44", x"22", 
    x"49", x"22", x"4F", x"22", x"55", x"22", x"5B", x"22", x"61", x"22", x"67", x"22", x"6D", x"22", x"72", x"22", 
    x"78", x"22", x"7E", x"22", x"84", x"22", x"8A", x"22", x"90", x"22", x"96", x"22", x"9B", x"22", x"A1", x"22", 
    x"A7", x"22", x"AD", x"22", x"B3", x"22", x"B9", x"22", x"BE", x"22", x"C4", x"22", x"CA", x"22", x"D0", x"22", 
    x"D6", x"22", x"DC", x"22", x"E2", x"22", x"E7", x"22", x"ED", x"22", x"F3", x"22", x"F9", x"22", x"FF", x"22", 
    x"05", x"23", x"0A", x"23", x"10", x"23", x"16", x"23", x"1C", x"23", x"22", x"23", x"28", x"23", x"2E", x"23", 
    x"33", x"23", x"39", x"23", x"3F", x"23", x"45", x"23", x"4B", x"23", x"51", x"23", x"56", x"23", x"5C", x"23", 
    x"62", x"23", x"68", x"23", x"6E", x"23", x"74", x"23", x"7A", x"23", x"7F", x"23", x"85", x"23", x"8B", x"23", 
    x"91", x"23", x"97", x"23", x"9D", x"23", x"A2", x"23", x"A8", x"23", x"AE", x"23", x"B4", x"23", x"BA", x"23", 
    x"C0", x"23", x"C6", x"23", x"CB", x"23", x"D1", x"23", x"D7", x"23", x"DD", x"23", x"E3", x"23", x"E9", x"23", 
    x"EF", x"23", x"F4", x"23", x"FA", x"23", x"00", x"24", x"06", x"24", x"0C", x"24", x"12", x"24", x"17", x"24", 
    x"1D", x"24", x"23", x"24", x"29", x"24", x"2F", x"24", x"35", x"24", x"3B", x"24", x"40", x"24", x"46", x"24", 
    x"4C", x"24", x"52", x"24", x"58", x"24", x"5E", x"24", x"63", x"24", x"69", x"24", x"6F", x"24", x"75", x"24", 
    x"7B", x"24", x"81", x"24", x"87", x"24", x"8C", x"24", x"92", x"24", x"98", x"24", x"9E", x"24", x"A4", x"24", 
    x"AA", x"24", x"AF", x"24", x"B5", x"24", x"BB", x"24", x"C1", x"24", x"C7", x"24", x"CD", x"24", x"D3", x"24", 
    x"D8", x"24", x"DE", x"24", x"E4", x"24", x"EA", x"24", x"F0", x"24", x"F6", x"24", x"FB", x"24", x"01", x"25", 
    x"07", x"25", x"0D", x"25", x"13", x"25", x"19", x"25", x"1F", x"25", x"24", x"25", x"2A", x"25", x"30", x"25", 
    x"36", x"25", x"3C", x"25", x"42", x"25", x"48", x"25", x"4D", x"25", x"53", x"25", x"59", x"25", x"5F", x"25", 
    x"65", x"25", x"6B", x"25", x"70", x"25", x"76", x"25", x"7C", x"25", x"82", x"25", x"88", x"25", x"8E", x"25", 
    x"94", x"25", x"99", x"25", x"9F", x"25", x"A5", x"25", x"AB", x"25", x"B1", x"25", x"B7", x"25", x"BC", x"25", 
    x"C2", x"25", x"C8", x"25", x"CE", x"25", x"D4", x"25", x"DA", x"25", x"E0", x"25", x"E5", x"25", x"EB", x"25", 
    x"F1", x"25", x"F7", x"25", x"FD", x"25", x"03", x"26", x"08", x"26", x"0E", x"26", x"14", x"26", x"1A", x"26", 
    x"20", x"26", x"26", x"26", x"2C", x"26", x"31", x"26", x"37", x"26", x"3D", x"26", x"43", x"26", x"49", x"26", 
    x"4F", x"26", x"55", x"26", x"5A", x"26", x"60", x"26", x"66", x"26", x"6C", x"26", x"72", x"26", x"78", x"26", 
    x"7D", x"26", x"83", x"26", x"89", x"26", x"8F", x"26", x"95", x"26", x"9B", x"26", x"A1", x"26", x"A6", x"26", 
    x"AC", x"26", x"B2", x"26", x"B8", x"26", x"BE", x"26", x"C4", x"26", x"C9", x"26", x"CF", x"26", x"D5", x"26", 
    x"DB", x"26", x"E1", x"26", x"E7", x"26", x"ED", x"26", x"F2", x"26", x"F8", x"26", x"FE", x"26", x"04", x"27", 
    x"0A", x"27", x"10", x"27", x"15", x"27", x"1B", x"27", x"21", x"27", x"27", x"27", x"2D", x"27", x"33", x"27", 
    x"39", x"27", x"3E", x"27", x"44", x"27", x"4A", x"27", x"50", x"27", x"56", x"27", x"5C", x"27", x"61", x"27", 
    x"67", x"27", x"6D", x"27", x"73", x"27", x"79", x"27", x"7F", x"27", x"85", x"27", x"8A", x"27", x"90", x"27", 
    x"96", x"27", x"9C", x"27", x"A2", x"27", x"A8", x"27", x"AE", x"27", x"B3", x"27", x"B9", x"27", x"BF", x"27", 
    x"C5", x"27", x"CB", x"27", x"D1", x"27", x"D6", x"27", x"DC", x"27", x"E2", x"27", x"E8", x"27", x"EE", x"27", 
    x"F4", x"27", x"FA", x"27", x"FF", x"27", x"05", x"28", x"0B", x"28", x"11", x"28", x"17", x"28", x"1D", x"28", 
    x"22", x"28", x"28", x"28", x"2E", x"28", x"34", x"28", x"3A", x"28", x"40", x"28", x"46", x"28", x"4B", x"28", 
    x"51", x"28", x"57", x"28", x"5D", x"28", x"63", x"28", x"69", x"28", x"6E", x"28", x"74", x"28", x"7A", x"28", 
    x"80", x"28", x"86", x"28", x"8C", x"28", x"92", x"28", x"97", x"28", x"9D", x"28", x"A3", x"28", x"A9", x"28", 
    x"AF", x"28", x"B5", x"28", x"BB", x"28", x"C0", x"28", x"C6", x"28", x"CC", x"28", x"D2", x"28", x"D8", x"28", 
    x"DE", x"28", x"E3", x"28", x"E9", x"28", x"EF", x"28", x"F5", x"28", x"FB", x"28", x"01", x"29", x"07", x"29", 
    x"0C", x"29", x"12", x"29", x"18", x"29", x"1E", x"29", x"24", x"29", x"2A", x"29", x"2F", x"29", x"35", x"29", 
    x"3B", x"29", x"41", x"29", x"47", x"29", x"4D", x"29", x"53", x"29", x"58", x"29", x"5E", x"29", x"64", x"29", 
    x"6A", x"29", x"70", x"29", x"76", x"29", x"7B", x"29", x"81", x"29", x"87", x"29", x"8D", x"29", x"93", x"29", 
    x"99", x"29", x"9F", x"29", x"A4", x"29", x"AA", x"29", x"B0", x"29", x"B6", x"29", x"BC", x"29", x"C2", x"29", 
    x"C7", x"29", x"CD", x"29", x"D3", x"29", x"D9", x"29", x"DF", x"29", x"E5", x"29", x"EB", x"29", x"F0", x"29", 
    x"F6", x"29", x"FC", x"29", x"02", x"2A", x"08", x"2A", x"0E", x"2A", x"14", x"2A", x"19", x"2A", x"1F", x"2A", 
    x"25", x"2A", x"2B", x"2A", x"31", x"2A", x"37", x"2A", x"3C", x"2A", x"42", x"2A", x"48", x"2A", x"4E", x"2A", 
    x"54", x"2A", x"5A", x"2A", x"60", x"2A", x"65", x"2A", x"6B", x"2A", x"71", x"2A", x"77", x"2A", x"7D", x"2A", 
    x"83", x"2A", x"88", x"2A", x"8E", x"2A", x"94", x"2A", x"9A", x"2A", x"A0", x"2A", x"A6", x"2A", x"AC", x"2A", 
    x"B1", x"2A", x"B7", x"2A", x"BD", x"2A", x"C3", x"2A", x"C9", x"2A", x"CF", x"2A", x"D4", x"2A", x"DA", x"2A", 
    x"E0", x"2A", x"E6", x"2A", x"EC", x"2A", x"F2", x"2A", x"F8", x"2A", x"FD", x"2A", x"03", x"2B", x"09", x"2B", 
    x"0F", x"2B", x"15", x"2B", x"1B", x"2B", x"20", x"2B", x"26", x"2B", x"2C", x"2B", x"32", x"2B", x"38", x"2B", 
    x"3E", x"2B", x"44", x"2B", x"49", x"2B", x"4F", x"2B", x"55", x"2B", x"5B", x"2B", x"61", x"2B", x"67", x"2B", 
    x"6D", x"2B", x"72", x"2B", x"78", x"2B", x"7E", x"2B", x"84", x"2B", x"8A", x"2B", x"90", x"2B", x"95", x"2B", 
    x"9B", x"2B", x"A1", x"2B", x"A7", x"2B", x"AD", x"2B", x"B3", x"2B", x"B9", x"2B", x"BE", x"2B", x"C4", x"2B", 
    x"CA", x"2B", x"D0", x"2B", x"D6", x"2B", x"DC", x"2B", x"E1", x"2B", x"E7", x"2B", x"ED", x"2B", x"F3", x"2B", 
    x"F9", x"2B", x"FF", x"2B", x"05", x"2C", x"0A", x"2C", x"10", x"2C", x"16", x"2C", x"1C", x"2C", x"22", x"2C", 
    x"28", x"2C", x"2D", x"2C", x"33", x"2C", x"39", x"2C", x"3F", x"2C", x"45", x"2C", x"4B", x"2C", x"51", x"2C", 
    x"56", x"2C", x"5C", x"2C", x"62", x"2C", x"68", x"2C", x"6E", x"2C", x"74", x"2C", x"7A", x"2C", x"7F", x"2C", 
    x"85", x"2C", x"8B", x"2C", x"91", x"2C", x"97", x"2C", x"9D", x"2C", x"A2", x"2C", x"A8", x"2C", x"AE", x"2C", 
    x"B4", x"2C", x"BA", x"2C", x"C0", x"2C", x"C6", x"2C", x"CB", x"2C", x"D1", x"2C", x"D7", x"2C", x"DD", x"2C", 
    x"E3", x"2C", x"E9", x"2C", x"EE", x"2C", x"F4", x"2C", x"FA", x"2C", x"00", x"2D", x"06", x"2D", x"0C", x"2D", 
    x"12", x"2D", x"17", x"2D", x"1D", x"2D", x"23", x"2D", x"29", x"2D", x"2F", x"2D", x"35", x"2D", x"3A", x"2D", 
    x"40", x"2D", x"46", x"2D", x"4C", x"2D", x"52", x"2D", x"58", x"2D", x"5E", x"2D", x"63", x"2D", x"69", x"2D", 
    x"6F", x"2D", x"75", x"2D", x"7B", x"2D", x"81", x"2D", x"86", x"2D", x"8C", x"2D", x"92", x"2D", x"98", x"2D", 
    x"9E", x"2D", x"A4", x"2D", x"AA", x"2D", x"AF", x"2D", x"B5", x"2D", x"BB", x"2D", x"C1", x"2D", x"C7", x"2D", 
    x"CD", x"2D", x"D3", x"2D", x"D8", x"2D", x"DE", x"2D", x"E4", x"2D", x"EA", x"2D", x"F0", x"2D", x"F6", x"2D", 
    x"FB", x"2D", x"01", x"2E", x"07", x"2E", x"0D", x"2E", x"13", x"2E", x"19", x"2E", x"1F", x"2E", x"24", x"2E", 
    x"2A", x"2E", x"30", x"2E", x"36", x"2E", x"3C", x"2E", x"42", x"2E", x"47", x"2E", x"4D", x"2E", x"53", x"2E", 
    x"59", x"2E", x"5F", x"2E", x"65", x"2E", x"6B", x"2E", x"70", x"2E", x"76", x"2E", x"7C", x"2E", x"82", x"2E", 
    x"88", x"2E", x"8E", x"2E", x"93", x"2E", x"99", x"2E", x"9F", x"2E", x"A5", x"2E", x"AB", x"2E", x"B1", x"2E", 
    x"B7", x"2E", x"BC", x"2E", x"C2", x"2E", x"C8", x"2E", x"CE", x"2E", x"D4", x"2E", x"DA", x"2E", x"E0", x"2E"
    );

  shared variable coef : mtype := coef_init;
  signal douta_reg, ram_data_a : unsigned(7 downto 0) := (others => '0');
  signal doutb_reg, ram_data_b : unsigned(7 downto 0) := (others => '0');
begin
  porta: process (clka, addra, dia, ena, wea) is

  begin  -- process porta
    if rising_edge(clka) then
      if ena = '1' then
        douta <= coef(to_integer(addra));
        if wea = '1' then
          coef(to_integer(addra)) := dia;
        end if;
      end if;
    end if;
  end process porta;

  -- douta_register: process (clka) is
  -- begin  -- process douta_register
  --   if rising_edge(clka) then
  --     if regcea = '1' then
  --       douta_reg <= ram_data_a;
  --     else
  --       douta_reg <= (others => 'Z');
  --     end if;
  --   end if;
  -- end process douta_register;

  -- douta <= douta_reg;
  
  portb: process (clkb, addrb, dib, enb, web) is
    
  begin  -- process portb
    if rising_edge(clkb) then
      if enb = '1' then
        doutb <= coef(to_integer(addrb));
        if web = '1' then
          coef(to_integer(addrb)) := dib;
        end if;
      end if;
    end if;
  end process portb;
end beh;
